    Mac OS X            	   2  �     �                                    ATTR;���  �   �  \                  �  \  %com.apple.metadata:kMDItemWhereFroms bplist00�_�https://attachment.fbsbx.com/file_download.php?id=364283610316987&eid=ASt3zhNNNcq0NH_g8RK90r4Eerk8E_reHbaPxnTGMM7Fo6cxqrrtHHdBjn5iWHW51Cc&ext=1347970406&hash=ASt3Q960LTm5cHI3_whttps://www.facebook.com/groups/281885715257497/286740474772021/?comment_id=286846648094737&notif_t=group_comment_reply   �                           6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           This resource fork intentionally left blank                                                                                                                                                                                                                            ��